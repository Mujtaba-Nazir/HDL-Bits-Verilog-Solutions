module top_module( output one );
	
	assign one = 1'b1;     // assigns 1 bit binary value equal to 1 to one.
	
endmodule